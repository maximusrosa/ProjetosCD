library verilog;
use verilog.vl_types.all;
entity mbr_mux8x1_8b_vlg_check_tst is
    port(
        Y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_mux8x1_8b_vlg_check_tst;
