library verilog;
use verilog.vl_types.all;
entity mbr_div_freq_1b_vlg_vec_tst is
end mbr_div_freq_1b_vlg_vec_tst;
