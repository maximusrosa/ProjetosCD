library verilog;
use verilog.vl_types.all;
entity mbr_decod3x8_vlg_sample_tst is
    port(
        e0              : in     vl_logic;
        e1              : in     vl_logic;
        e2              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end mbr_decod3x8_vlg_sample_tst;
