library verilog;
use verilog.vl_types.all;
entity mbr_teste_maj_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_teste_maj_vlg_check_tst;
