library verilog;
use verilog.vl_types.all;
entity mbr_teste_maj is
    port(
        s               : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic
    );
end mbr_teste_maj;
