library verilog;
use verilog.vl_types.all;
entity mbr_div_freq_5b_vlg_check_tst is
    port(
        Q               : in     vl_logic_vector(0 to 4);
        sampler_rx      : in     vl_logic
    );
end mbr_div_freq_5b_vlg_check_tst;
