library verilog;
use verilog.vl_types.all;
entity mbr_mux4x1_1b_vlg_check_tst is
    port(
        X               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_mux4x1_1b_vlg_check_tst;
