library verilog;
use verilog.vl_types.all;
entity mbr_teste_maj_vlg_vec_tst is
end mbr_teste_maj_vlg_vec_tst;
