library verilog;
use verilog.vl_types.all;
entity teste_mux8x1_vlg_check_tst is
    port(
        pin_name1       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end teste_mux8x1_vlg_check_tst;
