library verilog;
use verilog.vl_types.all;
entity mbr_mux2x1_8b_vlg_vec_tst is
end mbr_mux2x1_8b_vlg_vec_tst;
