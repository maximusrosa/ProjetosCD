library verilog;
use verilog.vl_types.all;
entity mbr_prova_vlg_vec_tst is
end mbr_prova_vlg_vec_tst;
