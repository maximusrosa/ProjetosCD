library verilog;
use verilog.vl_types.all;
entity mbr_bloco_arit_4b_vlg_vec_tst is
end mbr_bloco_arit_4b_vlg_vec_tst;
