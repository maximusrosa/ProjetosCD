library verilog;
use verilog.vl_types.all;
entity mbr_div_freq_1b_vlg_check_tst is
    port(
        D               : in     vl_logic;
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_div_freq_1b_vlg_check_tst;
