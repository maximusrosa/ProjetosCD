library verilog;
use verilog.vl_types.all;
entity mbr_circ1_vlg_check_tst is
    port(
        f1              : in     vl_logic;
        f2              : in     vl_logic;
        p1              : in     vl_logic;
        p2              : in     vl_logic;
        p3              : in     vl_logic;
        p4              : in     vl_logic;
        p5              : in     vl_logic;
        p6              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_circ1_vlg_check_tst;
