library verilog;
use verilog.vl_types.all;
entity mbr_reg_8b_vlg_vec_tst is
end mbr_reg_8b_vlg_vec_tst;
