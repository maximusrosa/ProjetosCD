library verilog;
use verilog.vl_types.all;
entity mbr_disp_7_seg_vlg_vec_tst is
end mbr_disp_7_seg_vlg_vec_tst;
