library verilog;
use verilog.vl_types.all;
entity mbr_disp_7_seg_vlg_check_tst is
    port(
        s6              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_disp_7_seg_vlg_check_tst;
