library verilog;
use verilog.vl_types.all;
entity teste_mux8x1_vlg_vec_tst is
end teste_mux8x1_vlg_vec_tst;
