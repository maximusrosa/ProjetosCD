library verilog;
use verilog.vl_types.all;
entity neander_vlg_vec_tst is
end neander_vlg_vec_tst;
