library verilog;
use verilog.vl_types.all;
entity mbr_div_freq_5b_vlg_vec_tst is
end mbr_div_freq_5b_vlg_vec_tst;
