library verilog;
use verilog.vl_types.all;
entity mbr_reg_1b_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mbr_reg_1b_vlg_check_tst;
