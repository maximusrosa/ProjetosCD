library verilog;
use verilog.vl_types.all;
entity mbr_cont_n_bits_vlg_vec_tst is
end mbr_cont_n_bits_vlg_vec_tst;
