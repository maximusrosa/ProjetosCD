library verilog;
use verilog.vl_types.all;
entity mbr_decod3x8_vlg_vec_tst is
end mbr_decod3x8_vlg_vec_tst;
