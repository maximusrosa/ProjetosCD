library verilog;
use verilog.vl_types.all;
entity mbr_mux4x1_1b_vlg_vec_tst is
end mbr_mux4x1_1b_vlg_vec_tst;
