library verilog;
use verilog.vl_types.all;
entity mbr_circ1 is
    port(
        f1              : out    vl_logic;
        p4              : out    vl_logic;
        p1              : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic;
        p2              : out    vl_logic;
        d               : in     vl_logic;
        c               : in     vl_logic;
        p5              : out    vl_logic;
        p3              : out    vl_logic;
        p6              : out    vl_logic;
        f2              : out    vl_logic
    );
end mbr_circ1;
