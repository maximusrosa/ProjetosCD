library verilog;
use verilog.vl_types.all;
entity mbr_mux8x1_8b_vlg_vec_tst is
end mbr_mux8x1_8b_vlg_vec_tst;
