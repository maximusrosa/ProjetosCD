library verilog;
use verilog.vl_types.all;
entity mbr_circ1_vlg_vec_tst is
end mbr_circ1_vlg_vec_tst;
